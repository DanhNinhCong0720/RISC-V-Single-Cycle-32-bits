library verilog;
use verilog.vl_types.all;
entity RISCV_SingleCycle_testbench is
end RISCV_SingleCycle_testbench;
